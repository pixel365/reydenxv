module model

pub struct PriceCategory {
	id int
	is_active bool
	name string
	description string
}
